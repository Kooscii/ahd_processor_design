library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use ieee.math_real.all;


entity tb_cpu is
--  Port ( );
end tb_cpu;

architecture Behavioral of tb_cpu is

    component cpu is
        Port ( clk : in std_logic;
               rst : in std_logic;
               sw : in std_logic_vector (15 downto 0);
               led : out std_logic_vector (15 downto 0);
               btn : in std_logic_vector (4 downto 0);
               -- 7-seg
               seg : out std_logic_vector (6 downto 0);
               an : out std_logic_vector (3 downto 0);
               dp : out std_logic;
               -- inst update
               prog_addr : in std_logic_vector (31 downto 0);
               prog_wd : in std_logic_vector (31 downto 0);
               prog_clk : in std_logic;
               -- debug signal
               debug_0 : out std_logic_vector (31 downto 0);
               debug_1 : out std_logic_vector (31 downto 0)
               );
    end component;
    
    signal clk : std_logic := '0';
    signal rst : std_logic;
    signal sw : std_logic_vector (15 downto 0);
    signal led : std_logic_vector (15 downto 0);
    signal btn : std_logic_vector (4 downto 0);
    -- 7-seg
    signal seg : std_logic_vector (6 downto 0);
    signal an : std_logic_vector (3 downto 0);
    signal dp : std_logic;
    -- inst update
    signal prog_addr : std_logic_vector (31 downto 0);
    signal prog_wd : std_logic_vector (31 downto 0);
    signal prog_clk : std_logic;
    -- debug signal
    signal debug_0 : std_logic_vector (31 downto 0);
    signal debug_1 : std_logic_vector (31 downto 0);
    
    constant clk_period : time := 10 ns;
    
    type PROG is array(0 to 511) of STD_LOGIC_VECTOR (31 downto 0);
    signal program : PROG := (
-- >>> start >>>
		x"00000011",
		x"10010001",
		x"1002ffff",
		x"14340010",
		x"16950001",
		x"16b60001",
		x"16d70001",
		x"16f80001",
		x"1019ffff",
		x"1b390010",
		x"101a001f",
		x"101bffff",
		x"1bfc0010",
		x"2c1cfffe",
		x"02ffe012",
		x"2efc0001",
		x"3000001a",
		x"02dfe012",
		x"2edc0001",
		x"3000002f",
		x"02bfe012",
		x"2ebc0001",
		x"3000000c",
		x"029fe012",
		x"2e9c0001",
		x"3000000c",
		x"100b1946",
		x"156b0010",
		x"0f2a5f91",
		x"016a5013",
		x"200a0032",
		x"100b51b2",
		x"156b0010",
		x"0f2a41be",
		x"016a5013",
		x"200a0033",
		x"100b01a5",
		x"156b0010",
		x"0f2a5563",
		x"016a5013",
		x"200a0034",
		x"100b91ce",
		x"156b0010",
		x"0f2aa910",
		x"016a5013",
		x"200a0035",
		x"3000005e",
		x"100beedb",
		x"156b0010",
		x"0f2aa521",
		x"016a5013",
		x"200a0036",
		x"100b6d8f",
		x"156b0010",
		x"0f2a4b15",
		x"016a5013",
		x"200a0037",
		x"3000000c",
		x"10030000",
		x"10040004",
		x"029fe012",
		x"2a9cfffe",
		x"029fe012",
		x"2e9cfffe",
		x"001f5813",
		x"156b0010",
		x"029fe012",
		x"2a9cfffe",
		x"029fe012",
		x"2e9cfffe",
		x"033f5012",
		x"016a5013",
		x"204a0032",
		x"04630001",
		x"2c83fff1",
		x"3000005e",
		x"10030000",
		x"10040002",
		x"029fe012",
		x"2a9cfffe",
		x"029fe012",
		x"2e9cfffe",
		x"001f5813",
		x"156b0010",
		x"029fe012",
		x"2a9cfffe",
		x"029fe012",
		x"2e9cfffe",
		x"033f5012",
		x"016a5013",
		x"204a0036",
		x"04630001",
		x"2c83fff1",
		x"3000000c",
		x"10030003",
		x"1c6a0032",
		x"206a001a",
		x"08630001",
		x"2443fffc",
		x"100bb7e1",
		x"156b0010",
		x"0f2a5163",
		x"016a4013",
		x"100b9e37",
		x"156b0010",
		x"0f2a79b9",
		x"016a4813",
		x"11070000",
		x"20430000",
		x"10030001",
		x"1004001a",
		x"00e93810",
		x"20670000",
		x"04630001",
		x"2464fffc",
		x"10030000",
		x"10040000",
		x"10050000",
		x"100d001a",
		x"100e0004",
		x"100f004e",
		x"1008001a",
		x"10090004",
		x"01094010",
		x"1c670000",
		x"00e83810",
		x"14eb0003",
		x"18ea001d",
		x"016a4013",
		x"20680000",
		x"01094810",
		x"1c87001a",
		x"00e93810",
		x"10060000",
		x"03498012",
		x"00075813",
		x"3000008b",
		x"156b0001",
		x"04c60001",
		x"24d0fffd",
		x"10100020",
		x"00075013",
		x"30000091",
		x"194a0001",
		x"04c60001",
		x"24d0fffd",
		x"016a4813",
		x"2089001a",
		x"04630001",
		x"04840001",
		x"246d0001",
		x"10030000",
		x"248e0001",
		x"10040000",
		x"04a50001",
		x"24afffdf",
		x"3000000c",
		x"1c0f0028",
		x"1c100029",
		x"1014001f",
		x"1c080000",
		x"01e87810",
		x"1c080001",
		x"02088010",
		x"10020001",
		x"1003000d",
		x"14440001",
		x"04850001",
		x"01f07012",
		x"01c07014",
		x"11cd0000",
		x"01d07012",
		x"01c07014",
		x"01af6812",
		x"01a06814",
		x"01ae4012",
		x"01004014",
		x"02903812",
		x"08ea0020",
		x"00084813",
		x"100b0000",
		x"28eb0003",
		x"15290001",
		x"056b0001",
		x"300000b5",
		x"100b0000",
		x"294b0003",
		x"19080001",
		x"096b0001",
		x"300000ba",
		x"01284813",
		x"1c880000",
		x"01097810",
		x"01f07012",
		x"01c07014",
		x"11cd0000",
		x"01d07012",
		x"01c07014",
		x"01af6812",
		x"01a06814",
		x"01ae4012",
		x"01004014",
		x"028f3812",
		x"08ea0020",
		x"00084813",
		x"100b0000",
		x"28eb0003",
		x"15290001",
		x"056b0001",
		x"300000ce",
		x"100b0000",
		x"294b0003",
		x"19080001",
		x"096b0001",
		x"300000d3",
		x"01284813",
		x"1ca80000",
		x"01098010",
		x"04420001",
		x"2443ffca",
		x"200f002a",
		x"2010002b",
		x"1c0f002a",
		x"1c10002b",
		x"1014001f",
		x"1002000c",
		x"14440001",
		x"04850001",
		x"1ca80000",
		x"02084011",
		x"028f3812",
		x"08ea0020",
		x"00084813",
		x"100b0000",
		x"28eb0003",
		x"19290001",
		x"056b0001",
		x"300000ea",
		x"100b0000",
		x"294b0003",
		x"15080001",
		x"096b0001",
		x"300000ef",
		x"01098013",
		x"01f07012",
		x"01c07014",
		x"11cd0000",
		x"01d07012",
		x"01c07014",
		x"01af6812",
		x"01a06814",
		x"01ae4012",
		x"01008014",
		x"1c880000",
		x"01e84011",
		x"02903812",
		x"08ea0020",
		x"00084813",
		x"100b0000",
		x"28eb0003",
		x"19290001",
		x"056b0001",
		x"30000103",
		x"100b0000",
		x"294b0003",
		x"15080001",
		x"096b0001",
		x"30000108",
		x"01097813",
		x"01f07012",
		x"01c07014",
		x"11cd0000",
		x"01d07012",
		x"01c07014",
		x"01af6812",
		x"01a06814",
		x"01ae4012",
		x"01007814",
		x"08420001",
		x"2c02ffca",
		x"1c080001",
		x"02088011",
		x"1c080000",
		x"01e87811",
		x"200f002c",
		x"2010002d",
		x"fc00011e",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff",
		x"ffffffff"
-- <<< end <<<
    );
    
begin

    clk <= not clk after clk_period/2;
    
    UUT_cpu : cpu
        port map (
            clk => clk,
            rst => rst,
            sw => sw,
            led => led,
            btn => btn,
            -- 7-seg
            seg => seg,
            an => an,
            dp => dp,
            -- inst update
            prog_addr => prog_addr,
            prog_wd => prog_wd,
            prog_clk => prog_clk,
            debug_0 => debug_0,
            debug_1 => debug_1);
    
    process
    begin
        
        -- reseting
        rst <= '1';
        sw <= (others => '0');
        btn <= (others => '0');
        prog_addr <= (others => '0');
        prog_wd <= (others => '0');
        prog_clk <= '0';
        wait for 200ns;
        
        -- 1000 cases
        for i in 1 to 1000 loop
            -- doing some changes in your program
            -- example:
            -- program(5) = x"12345678";
            
            -- programing
            rst <= '1';
            for k in 0 to 255 loop
                prog_addr <= std_logic_vector( TO_UNSIGNED(k*4, 32));
                prog_wd <= program(k);
                
                wait for clk_period/2;
                prog_clk <= '1';
                wait for clk_period/2;
                prog_clk <= '0';
            end loop;
            
            -- running
            rst <= '0';
            prog_addr <= std_logic_vector( TO_UNSIGNED(0, 32));
            wait;
            
            -- assert here 
            -- assert condition
            --    report message
            --        severity failure;
       end loop;
        
    end process;


end Behavioral;